
package req_ack_pkg;

 import uvm_pkg::*; 
 `include "uvm_macros.svh"
 `include "item_req_ack.svh"
 `include "sequencer_req_ack.svh"
 `include "driver_req_ack.svh"
 `include "driver_slv.svh"
 `include "monitor_req_ack.svh"
 `include "agent_req_ack.svh"
 `include "scoreboard_req_ack.svh"
 `include "environment_req_ack.svh"
 `include "sequence2_req_ack.svh"
 `include "sequence_slv.svh"
 `include "req_ack_test2.svh"
endpackage